module top_module ( 
    input p1a, p1b, p1c, p1d, p1e, p1f,
    output p1y,
    input p2a, p2b, p2c, p2d,
    output p2y );
    
    wire w1, w2, w3, w4;
    and a1(w1, p2a, p2b);
    and a2(w2, p2c, p2d);
    or o1(p2y, w1, w2);
    and a3(w3, p1a, p1b, p1c);
    and a4(w4, p1d, p1e, p1f);
    or o2(p1y, w3, w4);
endmodule