module top_module( 
    input a, 
    input b, 
    output out );
    and gate(out,a, b);
endmodule