module top_module( input in, output out );
    not gate(out, in);
endmodule