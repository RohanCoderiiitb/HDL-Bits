module top_module( 
    input a, 
    input b, 
    output out );
    nor gate(out, a, b);
endmodule