module top_module (
    input [4:0] a, b, c, d, e, f,
    output [7:0] w, x, y, z );
    wire[31:0] concat_vec;
    assign concat_vec = {a, b, c, d, e, f, 2'b11};
    assign w = concat_vec[31:24];
    assign x = concat_vec[23:16];
    assign y = concat_vec[15:8];
    assign z = concat_vec[7:0];
endmodule